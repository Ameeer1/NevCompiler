module main

fn main() {
	tokenize("hello world")
}
