module main

fn main() {
	println(tokenize("
fun main -> print(ln())
		"))
}
