module main

fn main() {
	println(tokenize("
fun main -> print(ln(60.76))
		"))
}
